/* Configuration AES */

`define ENCRYPT
//`define DECRYPT 
`define ROUND_3CLK
//`define ROUND_4CLK
`define ONE_KEY
//`define TWO_KEY_SWITCH
//`define TWO_KEY_AUTO