/* Configuration AES */

`define ENCRYPT
//`define DECRYPT 
//`define ONE_KEY
`define TWO_KEY